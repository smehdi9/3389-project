library ieee;
use ieee.std_logic_1164.all;
PACKAGE opcodes IS
   CONSTANT SUBA = 1;
   CONSTANT CMPA = 2;
   CONSTANT LDAI = 3;
   CONSTANT LDAD = 4;
   CONSTANT LDAX = 5;
   CONSTANT LDAF = 6;
   CONSTANT STAD = 7;
   CONSTANT STAX = 8;
   CONSTANT STAF = 9;
   CONSTANT JSR = 10;
   CONSTANT RTS = 11;
   CONSTANT LINK = 12;
   CONSTANT UNLINK = 13;
   CONSTANT BEQ = 14;
   CONSTANT BLT = 15;
   CONSTANT BLE = 16;
   CONSTANT BRA = 17;
   CONSTANT ADDA = 18;
   CONSTANT CLRA = 19;
   CONSTANT PUSHA = 20;
   CONSTANT PUSHX = 21;
   CONSTANT POPA = 22;
   CONSTANT POPX = 23;
   CONSTANT INCA = 24;
   CONSTANT DECA = 25;
   CONSTANT INCX = 26;
   CONSTANT DECX = 27;
   CONSTANT NOP = 0;
   CONSTANT SHRA = 28;
   CONSTANT SHLA = 29;
   CONSTANT HALT = 30;
END PACKAGE;
